LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TristateBuffer IS PORT (
  E : IN STD_LOGIC;
  D : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
  Y : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ENTITY;

ARCHITECTURE Behavioural OF TriStateBuffer IS
BEGIN
  PROCESS
  BEGIN
    IF (E = '1') THEN
    ELSE
      Y <= (OTHERS => 'Z');
    END IF;
  END PROCESS;
END ARCHITECTURE;
