ENTITY full_adder_2bit IS
END ENTITY;
