LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.UNSIGNED_STD.ALL;

ENTITY ALU IS PORT (
  clk : IN STD_LOGIC;
  sel : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
  A   : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
  B   : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
  F   : OUT STD_LOGIC_VECTOR (7 DOWNTO 0) := "00000000");
END ENTITY;

ARCHITECTURE Behavior OF ALU IS
BEGIN

END ARCHITECTURE;
