LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ParityChecker IS
  PORT (
    A : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    Y : OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE RTL OF ParityChecker IS
BEGIN
  PROCESS (A)
  BEGIN
    Y <= XOR A;
  END PROCESS;
END ARCHITECTURE;
