LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Accumulator IS PORT (
  clk : IN STD_LOGIC;
  rst : IN STD_LOGIC;
  we  : IN STD_LOGIC;
  Din : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
  Q   : OUT STD_LOGIC_VECTOR (7 DOWNTO 0));

END ENTITY;

ARCHITECTURE Behavioral OF Accumulator IS

BEGIN

END ARCHITECTURE;
